module full_adder(a, b, sum, carry);
endmodule