module top(); assign x = 1'b1; endmodule